/* verilator lint_off DECLFILENAME */
/* verilator lint_off UNUSED */
/*
    This is a testbench meant to test the cpu with a single port axi
    wrapper. The module contains an instantiation of a cpu that is 
    meant to be provided by the tester. 
    
    The device under test cpu must be named axi_cpu_wrapper. With an
    AXI4 single port. Our implmentation have additional buses that is
    not used for memory operation. These buses serve as a stopping point
    for the simulation. Read the simulation file for more information.

    Our modules are generated by Chisel. Hence the clock is named "clock".
    The reset is named "reset" and is an active high signal.
*/

module testbench ( 
    input        clock,
    input        reset,
    input        giveCtrlToCpu,
    output [7:0] storeOut_value,
    output       storeOut_valid,
    input        programmer_byteValid,
    input  [7:0] programmer_byte
);
    /*
        8 columns, 1023 rows
        column address is the last 3 bits of address
    */
    reg [7:0] mem [0:1023][0:7];

    reg [1:0]  AWID;
    reg [63:0] AWADDR;
    reg [7:0]  AWLEN;
    reg [2:0]  AWSIZE;
    reg [1:0]  AWBURST;
    reg        AWLOCK;
    reg [3:0]  AWCACHE;
    reg [2:0]  AWPROT;
    reg [3:0]  AWQOS;
    reg [3:0]  AWREGION;
    reg        AWVALID;

    reg [63:0] WDATA;
    reg [7:0]  WSTRB;
    reg        WLAST;
    reg        WVALID;

    reg  [1:0] BID;
    reg  [1:0] BRESP;
    reg        BVALID;

    reg [1:0]  ARID;
    reg [63:0] ARADDR;
    reg [7:0]  ARLEN;
    reg [2:0]  ARSIZE;
    reg [1:0]  ARBURST;
    reg        ARLOCK;
    reg [3:0]  ARCACHE;
    reg [2:0]  ARPROT;
    reg [3:0]  ARQOS;
    reg [3:0]  ARREGION;
    reg        ARVALID;

    reg [1:0]  RID;
    reg [63:0] RDATA;
    reg [1:0]  RRESP;
    reg        RLAST;
    reg        RVALID;

    wire [1:0]  temp_AWID;
    wire [63:0] temp_AWADDR;
    wire [7:0]  temp_AWLEN;
    wire [2:0]  temp_AWSIZE;
    wire [1:0]  temp_AWBURST;
    wire        temp_AWLOCK;
    wire [3:0]  temp_AWCACHE;
    wire [2:0]  temp_AWPROT;
    wire [3:0]  temp_AWQOS;
    wire [3:0]  temp_AWREGION;
    wire        temp_AWVALID;

    wire [63:0] temp_WDATA;
    wire [7:0]  temp_WSTRB;
    wire        temp_WLAST;
    wire        temp_WVALID;

    wire  [1:0] temp_BID;
    wire  [1:0] temp_BRESP;
    wire        temp_BREADY;

    wire [1:0]  temp_ARID;
    wire [63:0] temp_ARADDR;
    wire [7:0]  temp_ARLEN;
    wire [2:0]  temp_ARSIZE;
    wire [1:0]  temp_ARBURST;
    wire        temp_ARLOCK;
    wire [3:0]  temp_ARCACHE;
    wire [2:0]  temp_ARPROT;
    wire [3:0]  temp_ARQOS;
    wire [3:0]  temp_ARREGION;
    wire        temp_ARVALID;

    wire [1:0]  temp_RID;
    wire [63:0] temp_RDATA;
    wire [1:0]  temp_RRESP;
    wire        temp_RLAST;
    wire        temp_RREADY;

    reg [63:0] programAddress;
    wire [7:0] testResultData;
    
    axi_cpu_wrapper dutCore(
        .clock(clock),
        .reset(reset),

        .MEM_AWID(temp_AWID),
        .MEM_AWADDR(temp_AWADDR),
        .MEM_AWLEN(temp_AWLEN),
        .MEM_AWSIZE(temp_AWSIZE),
        .MEM_AWBURST(temp_AWBURST),
        .MEM_AWLOCK(temp_AWLOCK),
        .MEM_AWCACHE(temp_AWCACHE),
        .MEM_AWPROT(temp_AWPROT),
        .MEM_AWQOS(temp_AWQOS),
        .MEM_AWREGION(temp_AWREGION),
        .MEM_AWVALID(temp_AWVALID),
        .MEM_AWREADY(~AWVALID),

        .MEM_WDATA(temp_WDATA),
        .MEM_WSTRB(temp_WSTRB),
        .MEM_WLAST(temp_WLAST),
        .MEM_WVALID(temp_WVALID),
        .MEM_WREADY(~WVALID),

        .MEM_BID(BID), 
        .MEM_BRESP(2'b00), // all transaction will assumed to be complete
        .MEM_BVALID(BVALID),
        .MEM_BREADY(temp_BREADY),

        .MEM_ARID(temp_ARID),
        .MEM_ARADDR(temp_ARADDR),
        .MEM_ARLEN(temp_ARLEN),
        .MEM_ARSIZE(temp_ARSIZE),
        .MEM_ARBURST(temp_ARBURST),
        .MEM_ARLOCK(temp_ARLOCK),
        .MEM_ARCACHE(temp_ARCACHE),
        .MEM_ARPROT(temp_ARPROT),
        .MEM_ARQOS(temp_ARQOS),
        .MEM_ARREGION(temp_ARREGION),
        .MEM_ARVALID(temp_ARVALID),
        .MEM_ARREADY(~ARVALID),

        .MEM_RID(RID),
        .MEM_RDATA(RDATA),
        .MEM_RRESP(2'b00), // all transaction are assumed to be OKAY
        .MEM_RLAST(1'b1), // only supports burst length of 1
        .MEM_RVALID(RVALID),
        .MEM_RREADY(temp_RREADY),

        .giveCtrlToCpu(giveCtrlToCpu),
        .testResultData(testResultData)
    );
    assign storeOut_value = testResultData;
    assign storeOut_valid = 1'b0;
    always @(posedge clock) begin
        if (!AWVALID) begin
            // getting write address
            AWID        <= temp_AWID;
            AWADDR      <= temp_AWADDR;
            AWLEN       <= temp_AWLEN;
            AWSIZE      <= temp_AWSIZE;
            AWBURST     <= temp_AWBURST;
            AWLOCK      <= temp_AWLOCK;
            AWCACHE     <= temp_AWCACHE;
            AWPROT      <= temp_AWPROT;
            AWQOS       <= temp_AWQOS;
            AWREGION    <= temp_AWREGION;
            AWVALID     <= temp_AWVALID;
        end else if (WVALID && !BVALID) begin
            // data is available for write
            // one supports burst length on one
            // response buffer needs to be free
            AWVALID <= 1'b0; // operation completed within one cycle 
        end
        if (!WVALID) begin
            // getting write data
            WDATA <= temp_WDATA;
            WSTRB <= temp_WSTRB;
            WVALID <= temp_WVALID;
        end else if (AWVALID && !BVALID) begin
            // address is available for write
            // one supports burst length on one
            // response buffer needs to be free
            WVALID <= 1'b0; // operation completed within one cycle
        end

        if (AWVALID && WVALID && !BVALID && giveCtrlToCpu) begin
            // performing write
            // next buffer needs to be empty
            if (WSTRB[0]) mem[AWADDR[12:3]][0] <= WDATA[7:0];
            if (WSTRB[1]) mem[AWADDR[12:3]][1] <= WDATA[15:8];
            if (WSTRB[2]) mem[AWADDR[12:3]][2] <= WDATA[23:16];
            if (WSTRB[3]) mem[AWADDR[12:3]][3] <= WDATA[31:24];
            if (WSTRB[4]) mem[AWADDR[12:3]][4] <= WDATA[39:32];
            if (WSTRB[5]) mem[AWADDR[12:3]][5] <= WDATA[47:40];
            if (WSTRB[6]) mem[AWADDR[12:3]][6] <= WDATA[55:48];
            if (WSTRB[7]) mem[AWADDR[12:3]][7] <= WDATA[63:56];
        end else if (!giveCtrlToCpu && programmer_byteValid) begin
            mem[programAddress[12:3]][programAddress[2:0]] <= programmer_byte;
        end

        if (AWVALID && WVALID && !BVALID) begin
            BID <= AWID;
            AWVALID <= 1'b0;
            WVALID <= 1'b0;
            BVALID <= 1'b1;
        end else if (BVALID && temp_BREADY) begin
            BVALID <= 1'b0;
        end

        if (reset) begin
            programAddress <= 64'b0;
        end else if (programmer_byteValid && !giveCtrlToCpu) begin
            programAddress <= (programAddress + 64'b1);
        end

        if (!ARVALID) begin
            ARADDR      <= temp_ARADDR;
            ARVALID     <= temp_ARVALID;
            ARID        <= temp_ARID;
            ARLEN       <= temp_ARLEN;
            ARSIZE      <= temp_ARSIZE;
            ARBURST     <= temp_ARBURST;
            ARLOCK      <= temp_ARLOCK;
            ARCACHE     <= temp_ARCACHE;
            ARPROT      <= temp_ARPROT;
            ARQOS       <= temp_ARQOS;
            ARREGION    <= temp_ARREGION;
        end else if(!RVALID) begin
            // there is an request buffered
            ARVALID <= 1'b0;
            RID <= ARID;
            RVALID <= ARVALID;
            RDATA <= {
                mem[ARADDR[12:3]][7],
                mem[ARADDR[12:3]][6],
                mem[ARADDR[12:3]][5],
                mem[ARADDR[12:3]][4],
                mem[ARADDR[12:3]][3],
                mem[ARADDR[12:3]][2],
                mem[ARADDR[12:3]][1],
                mem[ARADDR[12:3]][0]};
        end

        if (RVALID && temp_RREADY) begin
            RVALID <= 1'b0;
        end

    end
endmodule